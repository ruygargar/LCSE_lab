--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   20:22:02 11/10/2013
-- Design Name:   
-- Module Name:   C:/Users/Silvia/Desktop/RS232 project/RS232/tb_RS232_TX.vhd
-- Project Name:  RS232
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: RS232_TX
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tb_RS232_TX IS
END tb_RS232_TX;
 
ARCHITECTURE behavior OF tb_RS232_TX IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT RS232_TX
    PORT(
         Clk : IN  std_logic;
         Reset : IN  std_logic;
         Start : IN  std_logic;
         Data : IN  std_logic_vector(7 downto 0);
         EOT : OUT  std_logic;
         TX : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal Clk : std_logic := '0';
   signal Reset : std_logic := '0';
   signal Start : std_logic := '0';
   signal Data : std_logic_vector(7 downto 0) := (others => '0');

 	--Outputs
   signal EOT : std_logic;
   signal TX : std_logic;

   -- Clock period definitions
   constant Clk_period : time := 50 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: RS232_TX PORT MAP (
          Clk => Clk,
          Reset => Reset,
          Start => Start,
          Data => Data,
          EOT => EOT,
          TX => TX
        );

   -- Clock process definitions
   Clk_process :process
   begin
		Clk <= '0';
		wait for Clk_period/2;
		Clk <= '1';
		wait for Clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      wait for 100 ns;	
      reset <= '1';
      wait for Clk_period*10;
		data <= "10101010";
		start <= '1';
		wait until EOT = '0';
		start <= '0';
		wait for 10 us;
		data <= "00000000";
		start <= '1';
		wait for 10 us;
		start <= '0';
		wait for 110 us;
		data <= "11001100";
		start <= '1';
		wait until EOT = '0';
		start <= '0';
      wait;
   end process;

END;
